VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO test
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 20 BY 10 ;
  SYMMETRY X Y R90 ;
  PIN avdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0 3.8 1.1 6 ;
    END
  END avdd
  PIN agnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 18.65 3.3 20 6 ;
    END
  END agnd
  PIN x
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 4.7 8.2 6.5 10 ;
    END
    PORT
      LAYER ME1 ;
        RECT 4.7 0 6.5 1.8 ;
    END
  END x
  OBS
    LAYER ME1 ;
      RECT 17.9 3.3 18.39 6 ;
      RECT 4.7 2.06 6.5 7.94 ;
      RECT 1.36 3.8 1.5 6 ;
    LAYER ME1 SPACING 0.16 ;
      RECT 6.82 6.32 20 10 ;
      RECT 0 6.32 4.38 10 ;
      RECT 1.42 2.12 18.33 7.88 ;
      RECT 0 0 4.38 3.48 ;
      RECT 6.82 0 20 2.98 ;
    LAYER ME2 SPACING 0.2 ;
      RECT 6.8 6.3 20 10 ;
      RECT 0 6.3 4.4 10 ;
      RECT 1.4 2.1 18.35 7.9 ;
      RECT 0 0 4.4 3.5 ;
      RECT 6.8 0 20 3 ;
    LAYER ME3 SPACING 0.2 ;
      RECT 0 0 20 10 ;
    LAYER ME4 SPACING 0.2 ;
      RECT 0 0 20 10 ;
    LAYER ME5 SPACING 0.2 ;
      RECT 0 0 20 10 ;
    LAYER ME6 SPACING 0.2 ;
      RECT 0 0 20 10 ;
    LAYER ME7 SPACING 0.4 ;
      RECT 0 0 20 10 ;
    LAYER ME8 SPACING 1.5 ;
      RECT 0 0 20 10 ;
  END
END test

END LIBRARY
